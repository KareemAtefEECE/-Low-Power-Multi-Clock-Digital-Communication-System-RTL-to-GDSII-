
module strt_check(
    input wire CLK,
    input wire RST,
    input wire sampled_bit,
    input wire enable,
    output reg strt_glitch
);

always @(posedge CLK, negedge RST) begin
    if(!RST) strt_glitch <= 1'b0;
    else if(enable) begin
        strt_glitch <= (sampled_bit != 1'b0)?1'b1:1'b0;
    end
end

endmodule